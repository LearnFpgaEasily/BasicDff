entity simple_dff is 
port (
    D   : in std_logic;
    CLK : in std_logic;
    RS  : in std_logic;
    CE  : in std_logic;
    Q   : out std_logic;
);
end entity;

architecture arch of simple_dff is

begin


end architecture;
